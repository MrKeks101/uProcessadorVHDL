library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port(
        clk       : in std_logic;
        address  : in unsigned(6 downto 0);
        data_out      : out unsigned(17 downto 0)
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(17 downto 0);
    constant conteudo_rom : mem := (
        0 => "00" & "0001" & "001" & "000100001",    
        1 => "00" & "0001" & "010" & "000000010",     
        2 => "00" & "0001" & "011" & "000000001", 

        3 => "00" & "0000000000000000", 
        4 => "00" & "0111" & "01" & "0000" & "010" & "010",  
        5 => "00" & "0011" & "010" & "011" & "000000", 
        6 => "00" & "0101" & "010" & "001" & "000000", 
        7 => "00" & "1101" & "11" & "000" & "0000100",      
        
        8 => "00" & "0000000000000000",
        9 => "00" & "0001" & "010" & "000000" & "100",
        10 => "00" & "0001" & "011" & "000000" & "010",
        11 => "00" & "0111" & "01" & "0000" & "010" & "000",
        12 => "00" & "0011" & "010" & "011" & "000000",
        13 => "00" & "0101" & "010" & "001" & "000000",
        14 => "00" & "1101" & "11" & "000" & "0001011",      
        
        15 => "00" & "0000000000000000",       
        16 => "00" & "0001" & "010" & "000000110", 
        17 => "00" & "0001" & "011" & "000000011", 
        18 => "00" & "0111" & "01" & "0000" & "010" & "000",  
        19 => "00" & "0011" & "010" & "011" & "000000", 
        20 => "00" & "0101" & "010" & "001" & "000000",     
        21 => "00" & "1101" & "11" & "000" & "0010010",      
        
        22 => "00" & "0000000000000000",       
        23 => "00" & "0001" & "010" & "000001010",       
        24 => "00" & "0001" & "011" & "000000101",      
        25 => "00" & "0111" & "01" & "0000" & "010" & "000",       
        26 => "00" & "0011" & "010" & "011" & "000000",
        27 => "00" & "0101" & "010" & "001" & "000000",      
        28 => "00" & "1101" & "11" & "000" & "0011001",     

        29 => "00" & "0000000000000000",     
        30 => "00" & "0001" & "001" & "000100000",     
        31 => "00" & "0001" & "010" & "000000010",         
        32 => "00" & "0001" & "011" & "000000001", 
        33 => "00" & "1000" & "100" & "010" & "000000", 
        34 => "00" & "0011" & "010" & "011" & "000000",
        35 => "00" & "0100" & "100" & "000" & "000000", 
        36 => "00" & "1101" & "10" & "000" & "0101000",
        37 => "00" & "0101" & "001" & "010" & "000000",  
        38 => "00" & "1101" & "11" & "000" & "1111111",
        39 => "00" & "1111" & "00000" & "0100001",
        40 => "00" & "0010" & "111" & "100" & "000000",
        41 => "00" & "1111" & "00000" & "0100001",
        others => (others=>'0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data_out <= conteudo_rom(to_integer(address));
        end if;
    end process;

end architecture;